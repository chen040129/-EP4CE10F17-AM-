library verilog;
use verilog.vl_types.all;
entity AM_vlg_vec_tst is
end AM_vlg_vec_tst;
